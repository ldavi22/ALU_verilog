module oddParityByte (
    input b0, b1, b2, b3, b4, b5, b6, b7,
    output p
);

assign p = ~ (b0 ^ b1 ^ b2 ^ b3 ^ b4 ^ b5 ^ b6 ^ b7);

endmodule

