module t_parityBit;


reg A,B,C;
wire D;

oddParityBitGenerator M1 (A,B,C,D);

initial
	begin
	A = 0; B = 0; C = 0;
	#20;
	A = 1; B = 0; C = 0;
	#20;
	A = 0; B = 1; C = 1;
	#20;
	A = 1; B = 0; C = 1;
	#20;

 $finish;
end
endmodule