module evenParityBitGenerator(A,B,C,D);

output D;
input A,B,C;

wire w1,w2,w3,w4,w5; 

not G1(w1,A);
xor G2(w2,B,C);
xnor G3(w3,B,C);
and G4(w4,w3,A);
and  G5(w5,w2,w1);
or G6(D,w5,w4);


endmodule